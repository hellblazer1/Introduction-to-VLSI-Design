* C:\Users\SAI ASHOK\q3_vlsi1.cir
G1 0 Vout N001 0 1000000
R1 Vin N001 1000
R2 Vout N001 3000
V1 0 Vin SINE(0 0.5 1000)
R3 Vout 0 1
.control
tran 50u 5m
run
*plot Vout Vin
wrdata plot1.dat Vout
wrdata plot2.dat Vin 
.endc
.end

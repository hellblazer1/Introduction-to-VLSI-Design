* C:\Users\SAI ASHOK\hw2_vlsi_q2.cir
.include "C:\Users\SAI ASHOK\TSMC180.lib"
.model nch_tt nmos
V1 n1 0 2.5
R1 n1 Vout 75k
C1 Vout 0 3p
M1 Vout Vin 0 0 nch_tt W=0.54u L=0.18u 
V2 Vin 0 PULSE(0 2.5 0 0 0 2u 4u)
.control
tran 0.01u 10u 6u
plot vout
meas tran OP max Vout
meas tran IP max Vin
let va = 0.1*OP
let vb = 0.9*OP
let vc = 0.5*IP
let vd = 0.5*OP
meas TRAN Tr TRIG V(Vout) VAL=va CROSS=1 TARG V(Vout) VAL=vb CROSS=1
meas TRAN Tf TRIG V(Vout) VAL=vb CROSS=2 TARG V(Vout) VAL=va CROSS=2
meas TRAN Tpl TRIG V(Vin) VAL=vc CROSS=1 TARG V(Vout) VAL=vd CROSS=1
meas TRAN Tph TRIG V(Vin) VAL=vc CROSS=2 TARG V(Vout) VAL=vd CROSS=2
print (tpl+tph)/2
.endc
.end
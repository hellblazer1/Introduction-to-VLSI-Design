* C:\Users\SAI ASHOK\q5_vlsi1.cir
V1 N001 0 PULSE(0 1 0 0.01n 0 5 5 0)
R1 Vout N001 1000
C1 Vout 0 0.000001
*control commands
.control
tran 0.1u 1ms
meas TRAN TIME_1 TRIG V(Vout) VAL=0 CROSS=1 TARG V(Vout) VAL=0.5 CROSS=1
plot vout
.endc
.end


